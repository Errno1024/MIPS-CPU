`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:22:55 11/07/2019 
// Design Name: 
// Module Name:    CTRL 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "def.v"
module CTRL(
	 input [31:0]instr,
	 input ben,
    output reg [`A3Slen-1:0] A3Sel,
    output reg [`WDSlen-1:0] WDSel,
    output reg [`SHSlen-1:0] SHSel,
    output reg [`ALUSlen-1:0] ALUSel,
    output reg [`NPCOp_len-1:0] NPCOp,
    output reg [`EXTOp_len-1:0] EXTOp,
    output reg [`ALUOp_len-1:0] ALUOp,
    output reg [`BJOp_len-1:0] BJOp,
	 output reg [`DMOp_len-1:0] DMOp,
	 output reg [`MDUOp_len-1:0] MDUOp,
    output RFWrB,
    output reg DMWr,
	 output reg MDUWr,
	 output reg[`TUselen-1:0] TUseRs,
	 output reg[`TUselen-1:0] TUseRt,
	 output reg[`TNewlen-1:0] TNew,
	 output reg `DMAS DMASel,
	 output reg `DMWS DMWSel,
	 output reg `TIndex TIndex,
	 output reg MDUDp, //MDU Dependence
	 output reg Likely,
	 output reg `EType EType,
	 output reg ILOP,
	 output reg eret,
	 output reg CP0Wr,
	 output reg jump
    );
	 reg RFWr,Bal,LinkUnconditionally;
	 assign RFWrB=
		( ~LinkUnconditionally & Bal ) ? ( RFWr & ben ) : RFWr;
	 
	 wire [5:0]opcode,funct;
	 wire [4:0]rs,rt,rd,shamt;
	 assign rs=instr[25:21],rt=instr[20:16],rd=instr[15:11],shamt=instr[10:6];
	 
	 assign opcode=instr[31:26],funct=instr[5:0];
	 wire[11:0]ins;
	 assign ins={opcode,funct};
	 wire[10:0]cop0;
	 assign cop0={rs,funct};
	 
always@(*)begin
	EType=`ET_NONE;
	ILOP=0;
	
	Bal=0;
	LinkUnconditionally=0;
	Likely=0;
	A3Sel=`A3S_rd;
	WDSel=`WDS_ALU;
	SHSel=`SHS_rs;
	ALUSel=`ALUS_rt;
	NPCOp=`NPC_PC4;
	EXTOp=`EXT_zero;
	ALUOp=`ALU_add;
	BJOp=`BJ_beq;
	DMOp=`DM_w;
	MDUOp=`MDU_lo;
	RFWr=0;
	DMWr=0;
	MDUWr=0;
	TUseRs=`TUse_N;
	TUseRt=`TUse_N;
	TNew=`TNew_E;
	DMASel=`DMAS_res;
	DMWSel=`DMWS_rt;
	TIndex=`TIndex_D;
	MDUDp=0;
	
	eret=0;
	CP0Wr=0;
	jump=0;
	casez(ins)
		`ins_addu:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_add;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_subu:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_sub;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_ori:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_or;
			EXTOp=`EXT_zero;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_lw:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_w;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_sw:begin
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_w;
			DMWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			
			EType=`ET_SAVE;
		end
		`ins_beq:begin
			NPCOp=`NPC_B;
			BJOp=`BJ_beq;
			TUseRs=`TUse_D;
			TUseRt=`TUse_D;
			jump=1;
		end
		`ins_lui:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_or;
			EXTOp=`EXT_high;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_j:begin
			NPCOp=`NPC_J;
			jump=1;
		end
		`ins_jal:begin
			A3Sel=`A3S_ra;
			WDSel=`WDS_NPC;
			NPCOp=`NPC_J;
			RFWr=1;
			TNew=`TNew_E;
			jump=1;
		end
		`ins_jr:begin
			NPCOp=`NPC_JR;
			TUseRs=`TUse_D;
			jump=1;
		end
		
		`ins_sll:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_sh;
			ALUSel=`ALUS_rt;
			EXTOp=`EXT_shift;
			ALUOp=`ALU_sll;
			RFWr=1;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
			if(instr==32'b0)begin//nop
				RFWr=0;
				TUseRs=`TUse_N;
				TUseRt=`TUse_N;
				TNew=`TNew_E;
			end
		end
		`ins_srl:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_sh;
			ALUSel=`ALUS_rt;
			EXTOp=`EXT_shift;
			RFWr=1;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
			ALUOp=`ALU_srl;
			case(rs)
				5'b00000:ALUOp=`ALU_srl;
				5'b00001:ALUOp=`ALU_rot;
			endcase
		end
		`ins_sra:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_sh;
			ALUSel=`ALUS_rt;
			EXTOp=`EXT_shift;
			ALUOp=`ALU_sra;
			RFWr=1;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_sllv:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_sll;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_srlv:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
			ALUOp=`ALU_srl;
			case(shamt)
				5'b00000:ALUOp=`ALU_srl;
				5'b00001:ALUOp=`ALU_rot;
			endcase
		end
		`ins_srav:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_sra;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_lh:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_h;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_lb:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_b;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_lhu:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_hu;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_lbu:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_bu;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_sh:begin
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_h;
			DMWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			
			EType=`ET_SAVE;
		end
		`ins_sb:begin
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_b;
			DMWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			
			EType=`ET_SAVE;
		end
		`ins_bne:begin
			NPCOp=`NPC_B;
			BJOp=`BJ_bne;
			TUseRs=`TUse_D;
			TUseRt=`TUse_D;
			jump=1;
		end
		`ins_jalr:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_NPC;
			NPCOp=`NPC_JR;
			RFWr=1;
			TUseRs=`TUse_D;
			TUseRt=`TUse_D;
			TNew=`TNew_E;
			jump=1;
		end
		`ins_slt:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_slt;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_sltu:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_sltu;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_slti:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_slt;
			EXTOp=`EXT_sign;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_sltiu:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_sltu;
			EXTOp=`EXT_sign;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_clo:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUOp=`ALU_clo;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_clz:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUOp=`ALU_clz;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_lwl:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_l;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_lwr:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_MEM;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_r;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			TNew=`TNew_W;
			
			EType=`ET_LOAD;
		end
		`ins_swl:begin
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_l;
			DMWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			
			EType=`ET_SAVE;
		end
		`ins_swr:begin
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			DMOp=`DM_r;
			DMWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_M;
			
			EType=`ET_SAVE;
		end
		`ins_bgtz:begin
			NPCOp=`NPC_B;
			BJOp=`BJ_bgtz;
			TUseRs=`TUse_D;
			jump=1;
		end
		`ins_blez:begin
			NPCOp=`NPC_B;
			BJOp=`BJ_blez;
			TUseRs=`TUse_D;
			jump=1;
		end
		`ins_ext:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_ext;
			EXTOp=`EXT_zero;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_ins:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_ins;
			EXTOp=`EXT_zero;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_movz:begin
			Bal=1;
			BJOp=`BJ_movz;
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_mov;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_D;
			TNew=`TNew_M;
		end
		`ins_movn:begin
			Bal=1;
			BJOp=`BJ_movn;
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_mov;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_D;
			TNew=`TNew_M;
		end
		
		`ins_mult:begin
			MDUOp=`MDU_mult;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end
		`ins_multu:begin
			MDUOp=`MDU_multu;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end
		`ins_mul:begin
			MDUOp=`MDU_mul;
			MDUWr=1;
			A3Sel=`A3S_rd;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end
		`ins_div:begin
			MDUOp=`MDU_div;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end
		`ins_divu:begin
			MDUOp=`MDU_divu;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end
		`ins_mfhi:begin
			MDUOp=`MDU_hi;
			MDUWr=0;
			A3Sel=`A3S_rd;
			WDSel=`WDS_MDU;
			RFWr=1;
			TNew=`TNew_M;
			MDUDp=1;
		end
		`ins_mflo:begin
			MDUOp=`MDU_lo;
			MDUWr=0;
			A3Sel=`A3S_rd;
			WDSel=`WDS_MDU;
			RFWr=1;
			TNew=`TNew_M;
			MDUDp=1;
		end
		`ins_mthi:begin
			MDUOp=`MDU_hi;
			MDUWr=1;
			TUseRs=`TUse_E;
			MDUDp=1;
		end
		`ins_mtlo:begin
			MDUOp=`MDU_lo;
			MDUWr=1;
			TUseRs=`TUse_E;
			MDUDp=1;
		end
		`ins_madd:begin
			MDUOp=`MDU_madd;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end		
		`ins_maddu:begin
			MDUOp=`MDU_maddu;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end		
		`ins_msub:begin
			MDUOp=`MDU_msub;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end		
		`ins_msubu:begin
			MDUOp=`MDU_msubu;
			MDUWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			MDUDp=1;
		end		
		
		`ins_add:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_add;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
			
			EType=`ET_ARIT;
		end
		`ins_sub:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_sub;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
			
			EType=`ET_ARIT;
		end
		`ins_and:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_and;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_or:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_or;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_xor:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_xor;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_nor:begin
			A3Sel=`A3S_rd;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_rt;
			ALUOp=`ALU_nor;
			RFWr=1;
			TUseRs=`TUse_E;
			TUseRt=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_addiu:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_addi:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_add;
			EXTOp=`EXT_sign;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
			
			EType=`ET_ARIT;
		end
		`ins_andi:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_and;
			EXTOp=`EXT_zero;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_xori:begin
			A3Sel=`A3S_rt;
			WDSel=`WDS_ALU;
			SHSel=`SHS_rs;
			ALUSel=`ALUS_imm;
			ALUOp=`ALU_xor;
			EXTOp=`EXT_zero;
			RFWr=1;
			TUseRs=`TUse_E;
			TNew=`TNew_M;
		end
		`ins_beql:begin
			Likely=1;
			NPCOp=`NPC_B;
			BJOp=`BJ_beq;
			TUseRs=`TUse_D;
			TUseRt=`TUse_D;
			jump=1;
		end
		`ins_bnel:begin
			Likely=1;
			NPCOp=`NPC_B;
			BJOp=`BJ_bne;
			TUseRs=`TUse_D;
			TUseRt=`TUse_D;
			jump=1;
		end
		`ins_bgtzl:begin
			Likely=1;
			NPCOp=`NPC_B;
			BJOp=`BJ_bgtz;
			TUseRs=`TUse_D;
			jump=1;
		end
		`ins_blezl:begin
			Likely=1;
			NPCOp=`NPC_B;
			BJOp=`BJ_blez;
			TUseRs=`TUse_D;
			jump=1;
		end
		
		`ins_bshfl:begin
			case(shamt)
				`bshfl_wsbh:begin
					A3Sel=`A3S_rd;
					WDSel=`WDS_ALU;
					ALUSel=`ALUS_rt;
					ALUOp=`ALU_wsbh;
					RFWr=1;
					TUseRt=`TUse_E;
					TNew=`TNew_M;
				end
				`bshfl_seb:begin
					A3Sel=`A3S_rd;
					WDSel=`WDS_ALU;
					ALUSel=`ALUS_rt;
					ALUOp=`ALU_seb;
					RFWr=1;
					TUseRt=`TUse_E;
					TNew=`TNew_M;
				end
				`bshfl_seh:begin
					A3Sel=`A3S_rd;
					WDSel=`WDS_ALU;
					ALUSel=`ALUS_rt;
					ALUOp=`ALU_seh;
					RFWr=1;
					TUseRt=`TUse_E;
					TNew=`TNew_M;
				end
			endcase
		end
		
		`ins_regimm:begin
			case(rt)
				`regimm_bgez:begin
					NPCOp=`NPC_B;
					BJOp=`BJ_bgez;
					TUseRs=`TUse_D;
					jump=1;
				end
				`regimm_bgezal:begin
					Bal=1;
					NPCOp=`NPC_B;
					BJOp=`BJ_bgez;
					A3Sel=`A3S_ra;
					WDSel=`WDS_NPC;
					RFWr=1;
					TUseRs=`TUse_D;
					TNew=`TNew_E;
					jump=1;
				end
				`regimm_bltz:begin
					NPCOp=`NPC_B;
					BJOp=`BJ_bltz;
					TUseRs=`TUse_D;
					jump=1;
				end
				`regimm_bltzal:begin
					Bal=1;
					NPCOp=`NPC_B;
					BJOp=`BJ_bltz;
					A3Sel=`A3S_ra;
					WDSel=`WDS_NPC;
					RFWr=1;
					TUseRs=`TUse_D;
					TNew=`TNew_E;
					jump=1;
				end
				`regimm_bgezl:begin
					Likely=1;
					NPCOp=`NPC_B;
					BJOp=`BJ_bgez;
					TUseRs=`TUse_D;
					jump=1;
				end
				`regimm_bgezall:begin
					Likely=1;
					Bal=1;
					NPCOp=`NPC_B;
					BJOp=`BJ_bgez;
					A3Sel=`A3S_ra;
					WDSel=`WDS_NPC;
					RFWr=1;
					TUseRs=`TUse_D;
					TNew=`TNew_E;
					jump=1;
				end
				`regimm_bltzl:begin
					Likely=1;
					NPCOp=`NPC_B;
					BJOp=`BJ_bltz;
					TUseRs=`TUse_D;
					jump=1;
				end
				`regimm_bltzall:begin
					Likely=1;
					Bal=1;
					NPCOp=`NPC_B;
					BJOp=`BJ_bltz;
					A3Sel=`A3S_ra;
					WDSel=`WDS_NPC;
					RFWr=1;
					TUseRs=`TUse_D;
					TNew=`TNew_E;
					jump=1;
				end
			endcase
		end
		`ins_cop0:begin
			casez(cop0)
				`cop0_mf:begin
					A3Sel=`A3S_rt;
					WDSel=`WDS_CP0;
					RFWr=1;
					TNew=`TNew_W;
				end
				`cop0_mt:begin
					CP0Wr=1;
					TUseRt=`TUse_M;
				end
				`cop0_eret:begin
					eret=1;
				end//eret should wait for mfc0 and mtc0!
			endcase
		end
		
		//Weird instructions
		
		//End of weird instructions
		default:begin
			ILOP=1;
		end
	endcase
end
endmodule
